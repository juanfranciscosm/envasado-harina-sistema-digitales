
module HOST_COM (
	probe,
	source);	

	input	[24:0]	probe;
	output	[16:0]	source;
endmodule
